module seven_seg_display
  (
    input clkIn,
    input rstIn);

endmodule